
/******************************
*** gen_fifo_defines_pkg    ***
*** Author: Ana Godoy       ***
*** Date: Jun 2024	    ***
*****************************/

package gen_fifo_defines_pkg;

  `define DATA_WIDTH    6'h20

endpackage
